`timescale 10ns / 10ps


module ScoreBoard
( 
    input   top_level_CLK50MHZ ,
    input  [1:0] top_level_KEY ,
    input  [3:0] top_level_SWITCH ,
    input  [12:0] top_level_DRAM_ADDR_i ,
    input  [15:0] top_level_DRAM_DATA_i ,
    input  [1:0] top_level_DRAM_BANK_ADDR_i ,
    input  [1:0] top_level_DRAM_DQM_i ,
    input   top_level_DRAM_RAS_N_i ,
    input   top_level_DRAM_CAS_N_i ,
    input   top_level_DRAM_CLK_EN_i ,
    input   top_level_DRAM_CLK_i ,
    input   top_level_DRAM_WR_EN_i ,
    input   top_level_DRAM_CS_N_i ,
    input   top_level_EEPROM_SCLK_i ,
    input   top_level_EEPROM_SDAT ,
    input   top_level_G_SENSOR_INT ,
    input   top_level_G_SENSOR_CS_i ,
    input   top_level_ADC_CS_N_i ,
    input   top_level_ADC_SADDR_i ,
    input   top_level_ADC_SDAT ,
    input   top_level_ADC_SCLK_i ,
    input   top_level_JP1_1 ,
    input   top_level_JP1_2_i ,
    input   top_level_JP1_3 ,
    input   top_level_JP1_4_i ,
    input   top_level_JP1_5_i ,
    input   top_level_JP1_6_i ,
    input   top_level_JP1_7_i ,
    input   top_level_JP1_8_i ,
    input   top_level_JP1_9_i ,
    input   top_level_JP1_10_i ,
    input   top_level_JP1_13_i ,
    input   top_level_JP1_14_i ,
    input   top_level_JP1_15_i ,
    input   top_level_JP1_16_i ,
    input   top_level_JP1_17_i ,
    input   top_level_JP1_18_i ,
    input   top_level_JP1_19_i ,
    input   top_level_JP1_20_i ,
    input   top_level_JP1_21_i ,
    input   top_level_JP1_22_i ,
    input   top_level_JP1_23_i ,
    input   top_level_JP1_24_i ,
    input   top_level_JP1_25_i ,
    input   top_level_JP1_26_i ,
    input   top_level_JP1_27_i ,
    input   top_level_JP1_28_i ,
    input   top_level_JP1_31_i ,
    input   top_level_JP1_32_i ,
    input   top_level_JP1_33_i ,
    input   top_level_JP1_34_i ,
    input   top_level_JP1_35_i ,
    input   top_level_JP1_36_i ,
    input   top_level_JP1_37_i ,
    input   top_level_JP1_38_i ,
    input   top_level_JP1_39_i ,
    input   top_level_JP1_40_i ,
    input   top_level_JP2_1 ,
    input   top_level_JP2_2_i ,
    input   top_level_JP2_3 ,
    input   top_level_JP2_4_i ,
    input   top_level_JP2_5_i ,
    input   top_level_JP2_6_i ,
    input   top_level_JP2_7_i ,
    input   top_level_JP2_8_i ,
    input   top_level_JP2_9_i ,
    input   top_level_JP2_10_i ,
    input   top_level_JP2_13_i ,
    input   top_level_JP2_14_i ,
    input   top_level_JP2_15_i ,
    input   top_level_JP2_16_i ,
    input   top_level_JP2_17_i ,
    input   top_level_JP2_18_i ,
    input   top_level_JP2_19_i ,
    input   top_level_JP2_20_i ,
    input   top_level_JP2_21_i ,
    input   top_level_JP2_22_i ,
    input   top_level_JP2_23_i ,
    input   top_level_JP2_24_i ,
    input   top_level_JP2_25_i ,
    input   top_level_JP2_26_i ,
    input   top_level_JP2_27_i ,
    input   top_level_JP2_28_i ,
    input   top_level_JP2_31_i ,
    input   top_level_JP2_32_i ,
    input   top_level_JP2_33_i ,
    input   top_level_JP2_34_i ,
    input   top_level_JP2_35_i ,
    input   top_level_JP2_36_i ,
    input   top_level_JP2_37_i ,
    input   top_level_JP2_38_i ,
    input   top_level_JP2_39_i ,
    input   top_level_JP2_40_i ,
    input   top_level_JP3_2 ,
    input   top_level_JP3_3 ,
    input   top_level_JP3_4 ,
    input   top_level_JP3_5_i ,
    input   top_level_JP3_6_i ,
    input   top_level_JP3_7_i ,
    input   top_level_JP3_8_i ,
    input   top_level_JP3_9_i ,
    input   top_level_JP3_10_i ,
    input   top_level_JP3_11_i ,
    input   top_level_JP3_12_i ,
    input   top_level_JP3_13_i ,
    input   top_level_JP3_15_i ,
    input   top_level_JP3_16_i ,
    input   top_level_JP3_17_i ,
    input reg [7:0] top_level_LED_i ,
    input   Stimulus_CLK50MHZ_o_i ,
    input  [1:0] Stimulus_KEY_o_i ,
    input  [3:0] Stimulus_SWITCH_o_i ,
    input  [12:0] Stimulus_DRAM_ADDR_i ,
    input  [15:0] Stimulus_DRAM_DATA_i ,
    input  [1:0] Stimulus_DRAM_BANK_ADDR_i ,
    input  [1:0] Stimulus_DRAM_DQM_i ,
    input   Stimulus_DRAM_RAS_N_i ,
    input   Stimulus_DRAM_CAS_N_i ,
    input   Stimulus_DRAM_CLK_EN_i ,
    input   Stimulus_DRAM_CLK_i ,
    input   Stimulus_DRAM_WR_EN_i ,
    input   Stimulus_DRAM_CS_N_i ,
    input   Stimulus_EEPROM_SCLK_i ,
    input   Stimulus_EEPROM_SDAT_o_i ,
    input   Stimulus_G_SENSOR_INT_o_i ,
    input   Stimulus_G_SENSOR_CS_i ,
    input   Stimulus_ADC_CS_N_i ,
    input   Stimulus_ADC_SADDR_i ,
    input   Stimulus_ADC_SDAT_o_i ,
    input   Stimulus_ADC_SCLK_i ,
    input   Stimulus_JP1_1_o_i ,
    input   Stimulus_JP1_2_i ,
    input   Stimulus_JP1_3_o_i ,
    input   Stimulus_JP1_4_i ,
    input   Stimulus_JP1_5_i ,
    input   Stimulus_JP1_6_i ,
    input   Stimulus_JP1_7_i ,
    input   Stimulus_JP1_8_i ,
    input   Stimulus_JP1_9_i ,
    input   Stimulus_JP1_10_i ,
    input   Stimulus_JP1_13_i ,
    input   Stimulus_JP1_14_i ,
    input   Stimulus_JP1_15_i ,
    input   Stimulus_JP1_16_i ,
    input   Stimulus_JP1_17_i ,
    input   Stimulus_JP1_18_i ,
    input   Stimulus_JP1_19_i ,
    input   Stimulus_JP1_20_i ,
    input   Stimulus_JP1_21_i ,
    input   Stimulus_JP1_22_i ,
    input   Stimulus_JP1_23_i ,
    input   Stimulus_JP1_24_i ,
    input   Stimulus_JP1_25_i ,
    input   Stimulus_JP1_26_i ,
    input   Stimulus_JP1_27_i ,
    input   Stimulus_JP1_28_i ,
    input   Stimulus_JP1_31_i ,
    input   Stimulus_JP1_32_i ,
    input   Stimulus_JP1_33_i ,
    input   Stimulus_JP1_34_i ,
    input   Stimulus_JP1_35_i ,
    input   Stimulus_JP1_36_i ,
    input   Stimulus_JP1_37_i ,
    input   Stimulus_JP1_38_i ,
    input   Stimulus_JP1_39_i ,
    input   Stimulus_JP1_40_i ,
    input   Stimulus_JP2_1_o_i ,
    input   Stimulus_JP2_2_i ,
    input   Stimulus_JP2_3_o_i ,
    input   Stimulus_JP2_4_i ,
    input   Stimulus_JP2_5_i ,
    input   Stimulus_JP2_6_i ,
    input   Stimulus_JP2_7_i ,
    input   Stimulus_JP2_8_i ,
    input   Stimulus_JP2_9_i ,
    input   Stimulus_JP2_10_i ,
    input   Stimulus_JP2_13_i ,
    input   Stimulus_JP2_14_i ,
    input   Stimulus_JP2_15_i ,
    input   Stimulus_JP2_16_i ,
    input   Stimulus_JP2_17_i ,
    input   Stimulus_JP2_18_i ,
    input   Stimulus_JP2_19_i ,
    input   Stimulus_JP2_20_i ,
    input   Stimulus_JP2_21_i ,
    input   Stimulus_JP2_22_i ,
    input   Stimulus_JP2_23_i ,
    input   Stimulus_JP2_24_i ,
    input   Stimulus_JP2_25_i ,
    input   Stimulus_JP2_26_i ,
    input   Stimulus_JP2_27_i ,
    input   Stimulus_JP2_28_i ,
    input   Stimulus_JP2_31_i ,
    input   Stimulus_JP2_32_i ,
    input   Stimulus_JP2_33_i ,
    input   Stimulus_JP2_34_i ,
    input   Stimulus_JP2_35_i ,
    input   Stimulus_JP2_36_i ,
    input   Stimulus_JP2_37_i ,
    input   Stimulus_JP2_38_i ,
    input   Stimulus_JP2_39_i ,
    input   Stimulus_JP2_40_i ,
    input   Stimulus_JP3_2_o_i ,
    input   Stimulus_JP3_3_o_i ,
    input   Stimulus_JP3_4_o_i ,
    input   Stimulus_JP3_5_i ,
    input   Stimulus_JP3_6_i ,
    input   Stimulus_JP3_7_i ,
    input   Stimulus_JP3_8_i ,
    input   Stimulus_JP3_9_i ,
    input   Stimulus_JP3_10_i ,
    input   Stimulus_JP3_11_i ,
    input   Stimulus_JP3_12_i ,
    input   Stimulus_JP3_13_i ,
    input   Stimulus_JP3_15_i ,
    input   Stimulus_JP3_16_i ,
    input   Stimulus_JP3_17_i ,
    input reg [7:0] Stimulus_LED_i 

);




endmodule
